package package_settings_v_6;
	parameter m1_6                                            = 16;
	parameter k_6															 = 13;
endpackage