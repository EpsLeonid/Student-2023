// ������ ��� ��������� ���� �����
module multiplier(

// ������� �����
input logic [7:0] A,
input logic [7:0] B,

// �������� ����
output logic [15:0] C

);

// ���������� �������� ��� �������� ����������
logic [15:0] result;

// ���� ������ �����������
always_comb begin

// �����������:
// ����� ���������� ���� ���������� - ��������� A �� B

// �������� A �� B
result = A * B;

// �����������:
// � ��������� ���������� �������� ��������� ���������

end

// �����������:
// �������� assign �������� �������� �� ����������� �������� result � ����� C

assign C = result;

endmodule