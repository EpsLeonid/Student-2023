module task_1(

//������ ������� ������
input wire [7:0] A,
input wire [7:0] B,
output wire [15:0] C
);
 assign C = A * B;  // ���������� ��������� � ������� ������ C// ���������� ��������� � ������� ������ C

endmodule