module zadanie_2 (
  input wire A,    // ���� A
  input wire B,    // ���� B
  output wire C    // ����� C
);

  assign C = A * B;  // ��������� �������� ��������� � ����������� ��������� ������ C

endmodule