module task1(

//������ ������� ������
input logic [7:0] A,
input logic [7:0] B,
output logic [15:0] C
);
 assign C = A * B;  // ���������� ��������� � ������� ������ C// ���������� ��������� � ������� ������ C

endmodule