import package_settings::*;
module reg8 (
	input wire [SIZE_A-1:0] A,
	input wire [SIZE_B-1:0] B,
	input wire [SIZE_C-1:0] C,
	input clk,
	//outputs
	output reg [SIZE_DATA_OUT-1:0] DATA_OUT );
	
	wire 	[SIZE_DATA_OUT-1:0] AB;
	assign AB[15:0] = A[7:0]*B[7:0]+C[7:0];
	

	
always @(clk)
	begin
		DATA_OUT[15:0] <= AB[15:0];
	end
endmodule