package package_settings_v_1;
	parameter M_1                                            = 16;
endpackage