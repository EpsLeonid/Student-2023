package package_settings_v_4;
	parameter M_4                                            = 16;
endpackage