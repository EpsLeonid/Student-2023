package package_settings_v2;
	//v2_filter-----------------------------------------------------------------
	parameter M_2                                            = 16;
	parameter k_2                                            = 5;
	parameter l_2                                            = 5;
	//--------------------------------------------------------------------------
endpackage