package package_settings;
//-----------------------------------------------------------------------------
	parameter SIZE_A                                  			= 8;
	parameter SIZE_B			                                 = 8;
	parameter SIZE_C		                                    = 16;
	parameter SIZE_DATA_OUT                                  = 17;
//-----------------------------------------------------------------------------
endpackage