package task_4;
	parameter SIZE_A                                  			= 8;
	parameter SIZE_B			                                 = 8;
	parameter SIZE_C		                                    = 8;
	parameter SIZE_DATA_OUT                                  = 16;
endpackage