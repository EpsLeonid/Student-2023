package package_settings_v_2;
	parameter M_2                                            = 16;
endpackage